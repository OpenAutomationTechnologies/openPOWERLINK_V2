// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G4IUz8pUICJG2yjTpwK2Y/dcmsVM0iTR/nAxmFYQc5veL9KFzw5nBNGZjp/Ox41u
0ftMM92cIYaNe5atKFwQK+GIwTLm834+7kfVpNucSUAYuTg6fF+E/u0mqtELTb35
/Rv7LHQ+UIAlYghmBJzPzyOeA5mQUZHfLmmxi4G2SAk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14512)
udVNCNRk6jnrUzOEGZ8dK2TcpAnaUtvl/erBFFr7xcFdPfNEQf82FmuWrvi8BrvZ
+AD7IqjdkLV7R7wEtL+yN98DVypvx+0Mu4u4EVKDKSoU9ogzageZPlmNCumpq+Jz
X8iZC9JJkvwB1EBOGk8va9yexLK9J4K8ly6XSNxmskdK0/5AI+eEPfEZF0qY1DXK
AVhYfxPInV8+opKoJy8WQGtrBamPB6E1Ikn8rt9htXMsH+OeaWmiSW+ZVqxVKO2E
cJHCKCErnE1QwkyROMry8hLYzMtYIsUgkm0vjZkzGzfTN0wGpwtbKv+Se4Uwl0dr
+hBHPLFKkKXTEeaSdO08aFc9FDtAX6ADQZtXYkQzhuD2zNdi4CBBG+IlYMlvjeyM
lTolvFhU9pIXL1K4udJm2eYX2EiOn0tErlWTSMUzNesSYV7BTdJHhT/TRt9Nnkst
DCX31uepn5uqmfZshgPe3z2V5pvCZwaTwvfSzDJ3IfYmujXmJp1XF//F6GrVyz79
FW4jY3M0AMgQmJYkbBOirUv1TzurIlWYlb/tDyHgXR7kgV/EFYpRFe1zrWqswf8L
ysyBvt/xwlMQYM5MsEid22LCmUkr7tprFWBXKcUcLCT+aTxkigsdRmrEoLZiKBFp
41cPbbkX/vgG2lo5yEPxDNpLcqbBqurhAmbqVoJJgjnb2xjqtDgkcjdFmuMDU4gz
7j2oE586yB5QLO6qOSKOAycg62orhuMA3ft8nrdhtS3/5uHfQRAtDdWT34lYz++E
jYDd+wdvDnB1x+mp48cqRPPiQuvnilhvsknXc5y8YoFUKySeDBMielpKD6X7gdTz
XiULoxg8wXvIPq0CFFjWBuYJMbNWm+gbqO7D54EHAP3RD8X4oIIQHOHznyJTKMHa
8raRohc+w7xGVnK8EmQ8/vUJbSOVWdABZelW4LbqPa8hAUnJaDZC95Noqp1dnUBx
FfQag082Tj2T5iJp2PisvrJgYRzshgzGU3ZsR0HUxHDTiVtT/aM3U5zO53AaURMX
owJ6MT/l2NeDpU+0sJ8aoUIzNJr0LhPlbb9+6xSwSPPgS8OVFHKVYcN4QYt8y/4Y
BgipwD4/L+KaCmxQqPKb53niaB83WPTTKBWZepQVSJLBGAzDWWgtTDq/FnVe51cl
Ud1Ch7woyoqKgVGpE03JXKFPV+o+is8HirmiFe+ePbTQ3afpxKa3NZzMgBm/wvkS
tXO9s96szSTD3QdE7DfCX1UpeDLOckJ3iQIYgb2HbBIBAIJXtSPqRuBAA03sBaep
bm3el7rt5tbWhZDqR/tordowr+VRG62IKdMSgXUsG8SaxQsnseqFd3BnVuZnFNia
cmcKHhSDqJ6IdN996Rn3iaCQmtlkHRJQ0QKNzkSlZ1G9FSNuCQULlD+ym+9qfAX/
OAtmUFRXs4KoD02uJtDxtIz1yVHIrN7stXHmvOAMy+CrdLQEScVQxV9jJ0RK9URa
4fAj+PVsGh3rJpWK9E8bXu/6y5i8HUqV172STs+KtuwMHbG2w4lCcLuGB3CE3lfr
pjrC6K3ZPkKATG6O+1dtzqY9ouBC5WkrV0S/yohxoFn1+xO3ubaNwaPsZej8y0J0
giNZ2CZdau6008uwYjo+qYPYuQKZ0nTvbbJcsps+8tvGInzpsTGnn7ueyOPCOlbB
IBt6dMRvLL7vpvfn7LnTg3PzdHgdifzEtgmiDmK8LSn23ZzSzh2ZPuL8tbNXMy7x
A82Eg6Ca9nrugHRzpNmXt82aamU3JraL5Tzc9nW5/wKMdI9EwYSzNIMWBoHr5arQ
PBN6dnsx7ZMq8K0qXJ+e77n/roFctQtoA1l4KRShXb2/zjhliFiBrswn8MFDPKSF
XzrCBmiu6uyNuQfHr+BgAoMlmuWpEZ5+k7se2Wrq8YEls5FadG2KBHOrw0gVd1Qn
ICX+orJ+IJW9iRiB5OMdaY3WZzgb3U7FXfNgBgn/grGo+8eVEjvFEd+I/HA1C8NP
eAQ8EHYNqsH+ghFQPw4tp5xAANfxVWAMlHu0h79cwSVjYBeo1BPecxhdgeyfCofs
cV6n47Al6HJ/Vf0yYzMPk51RTxMIkMH0mll4N/XbHKnP/cjAljLewVZeuhVsUanu
xqe07VvoQS7QV+BX99+w0fMF2+Ea2Fi7C/9l35QFA85Y5oA8WmyVK7AEDEnbCL4Z
CZAJrhFrST92eMEOWwRFOmc/f4UeC/0d01za7jMXabV3XAndKLvKC+LCbYxhGBfx
G7IuhRHP7lqTp/BTJnxogr1F/Nv94LL0rrMwPVbNflfNPPhswiX2W4DijM3uSl92
nvnms+zU7DGR7s+poHf2e6UyNPaK4fRPuPLGie6XImKGK6WoUAbQoQ2S97Ux35Ph
D+nVyp+eDFvJv0GsfyhUsR0mYFglfq7KRS/AoZ4hdSl3+F3Biitrwsr8EX2+FuVk
ct0unlkoD7NZD3fj3d2BXkELnG4PVe8hKEHYZPogi3qHEIJnrlp+JrBA5QbhMqZ/
q7Eqsu2H3VC2UjUPZ5BYKfjNMwKBBmvqPBtgEuuG/2l0WpDbTXay6I67FxNX4SHN
mIUZpFCDtsENZCmIBUCPAhsyYq6RzqSFwynCwzFvFWd3nva/nXpF1GC9vSInAypp
D2mIJt03ERWpFx90I/3vMnOlfcsjB+sLGrPpEEkuImFS5lhTywgBMHyLuUm0lZSF
cf/5tw82bq/gYXl3CVZesNAGaGnGKZdSSbjWG/J/ALfqjqf0MZMnn2IZjNcFzDqh
iIp2mkbPMyI7RkvASel8sNKXRiVGm6qZwE6Kq94ztLHXsuXz2gyNlqSai75rNUNJ
K1c4Q+1NcrJLgwFro3o7s2UGJ6UdGCO7XtUzEJG2x+grcoy6yebk7ybSpNUO33XA
7fzZHbrl/H9qyXSg/2EZv5oD4tiNO3BeGPw1+rEg4dyyg3yFYY+Y0iSEMT9+RHoo
3P9efFOcNjSkOPpCxB1V8sB/05/CCcOGTCBZcolUcPuhziTO8zFoc6BNAwyIkAtA
cCU1hshsq/Upq1AZSOoBaa6MbAecfxvvrAqV2RD1Vd8e/bCLIZhN3oehUAUQ7rRy
a19ihrtuAWla/nz/Ba3WwLt3oWhR8s9gnVg56qJ0H3qZrMJT34xuxveWrLrLaSmi
AdQRRNGPPve6gxvSDRMek7T2ElYtlLaeG602m1si40YyTWLxIsXLA7F8Jt5mVQRo
BKw4LCwKjfZsB3E6ehW8TgI5IUAsJvxrtwkFGDvhdjGYpJn5bGmYPPjTrq5bt2Wa
fVXKkI19V5Dvj3JDU9CiM5zT315C2tsdrae16N79wRGCI6TJksgtkXc8CJzbUkuL
cPpY0A8XSd5o8jGthEn9cvDOt08ORZI7uwAXZmMa6Ht19QgXoMueSezifCg58tbm
urWiqbJy8pujmW9KOJZjyu8lQgd1Bu6AtslZIBw1L1cU7FARci6PktRf0DJ0Dg6O
aRnGa84Sm7VhOmjRTboOScVSvjHmL5/wMdhuWJwVxCDitU2gbnEWRmGwcFJN8ty8
iivg09uhSrV53Oe82HSj8FIW3j9uSGePQDfKa1vCQC/pcHGhVsk8u/rlJknnGMCg
2EUa1KtjtLv3YF9TMw7EKbcL5Bii0+RLLdtOxK8L+71XF9L+hQ1Q4HhE4kB94LY9
/CCSRiDCnhXimYx404tUtE10SPfVU0g4ompySGNEsJHNsijt0qgnA7KhTPJLVyCA
3ccr5o//Zf21UA0TZZc3cNnRFN1aP0DN2cZCl3YJQqSWUNDfsInlHePm+LFLeBYD
uhinhe9JNgoaRe3TOGVRqCH9oVVofLBIsd9tBrV3ltuftWUPB/n+bUcX3MvP7c+y
aCWs16jUfOCW3LLLuju7zAA+fz7gxoCGf6qWX6jyVw7FHlOsIimMrLHcGGrzuF6W
2l5xG0ua1XBxJKqNABjUIeKHog+s26hK9aToHgXkMnotPAPF5WRmZxHlxR23B13t
mTQeBlHmmmVQmArVKTUnJo2pG7SyCKKH6jslA6BDBK4y8qYdnVPhVne8F1mpPQ/s
N9ihR+dVbsJoEBNL7xI7ssXIvLdPaF9TDgvIuNDJYby1HWvyN+VXjdmvvk9wEB+i
XbyRHj4fzds0o54tlzitOGwiQeZTzq97kgRgEzZSEoRYbcs47nrXOqC4ae3g1d/U
H6HJ0vK6eVOaMYPrCi4UeQsGuqdWgUGCKznC+VSZrjTS+O6EM8+EqdtqrVIud0K2
HXWXbFGro1vwZJMCKPDaYA+cwN16ycc1Rbe7z/SblTwKmnIvrJ4dn1xf0FktQxte
xMCmyU2cFz/vxLSboCSP/XLWnz8tCsIIKDmXWAGxAhRjkSbAIHNN1lm0YoJLLu4q
CODARLhOtDj4HjwS4HGvk8AC7RzFxtRCxUtLEFRPdM1nrhIN9+09NbTzBMyG7aRe
gsIU1Ovt76rf7U4GowQsQi+ve+yWMWTpE33aN70cSEElY/+nWrb4PHO4ZWRCF9KY
23P1PmhBsK+Q0M2Nx9DhcAVsK5Ljr9oeaCaZLP4yUlRlhnYPzup5yf/U+ienlJLV
FtGjCYgMW0/HSaB5LzRvgvlU+datHCqLoN8Tc8ijNi2pGSZpkcJ2hmgX0MauIEhd
Grj8oeFVYPjdpDmkGYETlsl8HmAao1PyQjvpvgU1DXsSqLvr6nmK/j391dw3TxKp
NtpIp053AsvdSYvA7lR2GnKtqFQgPfSk29aNTK74ZECJHqka9TGXjO0P2EDA8Mvu
PUZamlsgDyxTey5AB90t5SqVmgtB7wo5TsPV3UMR+vFJjpoJniZN30ckCxYINW/v
Z5xpN3j3+mNf/wZMnm/LSRqb458vuz+gv/J+w1+uXu30/IyYqchVktuERKh/rZp9
QgYgB32EOCXBg6iNAItuga9wzMQQdLOt32gGgFAQSdN65808QwBm1YNVu64iaCRu
KT4QybdMTTzLqK4ADi5eD13rZUiIpvPTYbfGPrq7Q5/KL0WwPzi+52Zsh8ypuox1
GrgZoaCKAW6kqGtGHTj20IcrpbrlgXDFv+nYVU78xduZocgaKGxI9Osdjby6DmlW
MWQWo9TYB24LCarlU6KYmBBXv0ZwQ7lNdGLKMDYAqIP+kritEGvI/KhdQn3ON7kJ
miVDx2KFJRop1QhxjZZlPtrz0mDZIDWBf4WmewprAldVR0RUior89CH5+ZGcQSLD
BLQ1stKYA+0O2dsHpxOQiFcYRkGjNRjuJYzik6fTcBV7zcs2ybL3Mu0n6ubB5mbi
Z6ZBoKuHqpZoYSQQE/h9AgC1SQniau/Z1boB6hn3Mj/dKzDzdvx6GZoY/whYmjKe
/dRv1ElzUw1996oPLAd8vbt9UmZshbAvZp+FMC6giI786QiYAzKfhjiGufEmydbC
l5ckPvWZu9/OhIztO4g0cqitxkKtO+IWAN2Xif8z9hyvwScMVIAk4NaIPafLSpIE
YdUOEZc59dKn5J9Y1Qruy1g9PbrskVQl3Rr9MsH6dVBpPUEXLTohVyOYUZzowMFs
8+itQrsafH8ZWNvjSop6CfCJz+umBqVfChcPI2+xot/3jNi3aE8TuHWAbHC9+JT4
SnwsyOy/gMjTGL5j9Vl2QIyF9Nc6e0wINwZcQ9ayhWNaDj509dCHXnfZJAyRYsNA
WgsIm20I+2NNpjkfaBJ+7hirKGYMmHvV8b5VGv1JE7TVBGmjTUUvN2BJD4GA2fuM
gkOVOgrUU7jbLXq9N7W1z8CsTEZtnaji/92HycnSaUPDl11rO+iZ2K0NML+QYZ3J
yAyyyzpQYNlni84Nn6TQpzPlIFGcfSwEDfk67kjT1BqsuQqKv/GwP4yr86W59zP5
5eSM37WEYeJLTpSpp/7LPSux+wqDoHOjGeD0wUc8P0tEDHSr8K8mnJjAUqI3CtBs
HPd+xlG5q+08Qaqyz7OpIUpxHTb6//1KtKv+SICt0JfMARFKryYjJQ1t4sYFEPIx
y0/MWZLeT+mQQlvSFwI9YpxULqBMXCqMIaueRIxRt7ki2RdqL49h7QYAK24M67OC
0YsgpBdUzSOGkVIhu8qILFDAp5NYIymnchKg/jXbk7jG8Ofq4z76oXk7xO7/lc58
BMhN+pgYgIqunUH9PLIujreddRfb/Tpk+q9hou7mR+ExK9ptYyHcPd1YZeyAyUHX
6OEsq8b/9/U/GMgafrKutIdUzDb7t3LhnkfrsyCcNY8cJYnEKSfgnELsWLruSzhh
MG/pvCxcup1qlP5ljvsoe1XFx1q03hh4Zt2gwfxiLtizAHmD1vSrdxtjpu7RyriQ
4vUd52DREfoF8Z3SbKMKe9HqvEr+DYf+rgaW8hP7AZJNdPDnKTs5msZf5FNhlV3u
stTDsNL/rY59ccNl6YF1P/e5Wb057B3Cpdhw5AYtdSt2BUf5ynPguyXcXnprkDfX
gowSX15N9bD8YZcblct8HVK8bL64kv7uVEavOfu7OUqIBwh/BYAPGaYNa2Kc6w4G
3Ja3jW4v31So5J0VrNVCMx4uNFBJPJGqyohdtphmwdjy9oEU/jyB2ABRaWWZrIQd
vimpGBX2h1gfyHJnaUoVn3sN/Pvgg+f6N/4u987QwixRs/rXp/vmQaoiIVCy9c/w
ZqqmnaR4GfqaU7LU+Kn2KqVV0rUQlhD0Ik+8lGAme/A7MmW1n9ftFbZutaxB2Zj5
RHg5ASqsUbEoITCi2OENdm8ndzDa9xBVFJqFq8cOD1U9/ZvJ++0nDualePsKvxIZ
Av4HGa2rdN7/LhETcn9hSgXhOoFTTl4fSydrmcvHP43N6Cnon4FP+x3vCPxQyQHs
MveZPrTRq2rc8xq1bFUKc3WqlSJXqYiKGles1E2VeQSCgSdfM7UJLhMne8mnTYMq
CxKFcwnNrbFUQH1oJLTEzVVsjEo8K7GEnAK76sjntwuTkL+itBKDAAdu7hpFg0PE
O8TPfLfLAr3Oh8Y9m5A0F0JFygYOkwXT2baKv9vAgyhu2YuntqB1NFBllM+G1g4y
UwIBQOII2MVYXjoK/l04WtIB0MmpiVDFqzjWvY/uvwGoQkvR1UQS2SELOA0YROYj
qD7+94casRbw/C9SZJKhVQ6eQtIGHhYHXzen8v2m9mb5OHNt3rD/oPhUOtWESTC3
ZTRCa2rQqPYoFbLtAMSWSUASbCGpb0xYorqYtYjelGyzdPXbHP7m2hyAGpB8e8+f
ZaF7MajHCw1sdliHkBm5T+8K4IY2DhDJRtiJFvWCP6EVMvaK6Lv9z+IeFQuVS32N
MHvYSTNh0iIJKnc/PfAcqNGfZeIWhqpt8IvseICcfD2QXN4VprIwOU1xedWtXSme
ZY/pS9R8bVGPh5BF/CU7XW8DAedOPWJjUjISuRlPjFUTkwgVvC8Y1XExSwDJ3iuS
wzyBdihlZKFofledOlEFLx0GQ0WyiNCUFuXXlEPp0S6RckHvQ714TVhI8bsI5/+4
0XpRJy5fW+ZFFoSgVPK9TKtLh9hZPLCekBXWUPfvbaj0cL1i58P4naV+pmjC8DIQ
js4mcfnZh/sTSiSXDHCqD5wXzQdSUADmxLyDfXB7RZmztSTWKqDDIkqOunoWlwAX
a06TUF5pQ8jA0JGB+nwAGVaFUy230p3ag3RGMrwayd9XHoL8uryu0JkV4Pzxdb5D
Rnfo+i7WS8btmZqyB5AhzTnH+1knUbApFUwEbQ9QjebGb/lrseBDdOkEQWesBRjc
3GAjClqVY0MoMjjnsK/6PK33I3S9iXpcmrM3lx7ojKfusKBS9e1W78rrG19KtYYP
etNRHyHJQDr3oKRAHy/HQBpN1kxUF5+OAEfp/qhnNI4o7sdO73vBVeWMmue3PiSo
d5HBVHBPjz89BOnHtTC41cQGiGjFjRlp9uY2NjecZsu0BQQWfu4hky6ziMLunPrO
x4HPU1pF/2kqjsDZWyUECYl2WDAQOwndhuIsy6rgmMeUpIQvM0DtKDVpAdHdu58i
2TXwXuHUs11rFDVFEllVN/CBWakQhvm/C0riaT5gqB1+iq3dWTpi99/Ji/DxFrCr
oOHaQaAqWnI+eLAGc/zKM34CRiZgs4EI0Xf6b3jW8eDxvJhF2pQTRJbGs/wggYz7
jbfot/4M4gPTvMdl1pMx5wyJOsZlZLfiZXfn1QdLXACI5du6hi7Jfku5jtpnwITs
wnTh4esymRxvF7OZ2PKRBlZnD5iyUMnedskDpkogaFrPV+iekunHbJPOqHqEFILY
096mmet7jJiV0uXWJmpu2eiv7CNygbKY8gl3sWn+dtyePyuQN6e/JZc7eNI0AznG
ayq9uqKukMN7jdef0bqKpv+0Wev/19YYV5Vb2WlvFNbc4srXb3qdtKge9Obdf6ll
llHubdGgJbeplSy/XJf0KpVapIq3AYQmxGwCY1aLuZCqOYWeWEXKMIxVT/9Yml9P
DaxzgO0avQ75N/0hmgBX9Qry71+2hIPQJMCbW2+MhhZUCbVdSjeNuZ1+6Y2Q8Nmp
q6j0g0ushM4hioT5VbfTQsVztBMUqkhH5M6ZUvv25Xavy6tIUlFp94uekWhjJB6i
p8HmQBdp0CQmepSMLd1lcArZl2FaYuFynCZ6jCVIEgcHAZ1fASDJwF9egS5gZcun
kH8d6w4Ujzjr6+9bytkKvNdSF18Cm6mj66I2SjOv/dWC8gTiNmKuOTUFs0UKWw2L
HusZ9nbJJs6arsQda//0UeV2SigaC031X2lUMtHT3FuGoUJYIqPShutqRB0MI0Xd
pqHs0aO8nkmgZWWLuv+cl3FQMXAB7zUYfIRlsdmy8b4t07aLacpn0R1kVwWzQtLr
3VFAFKr7O4gFmszBLZ3Hj60tTi5t3O9PrT7GWeKTZb7vDUHEssYOjM1tHGXME0Ib
rn+Yiz20c+OsYhhBbueI75w3aRTWBmOeQiuveBDa3v0N08JFaTK8dnqvZVwhnyFn
o5/WZKLp4vNdhY+lPEiUl9rl6vClEsFDFBPIqs72q2muXdMkO1exAfKPIIzv2iWB
5ua1vlTd28VrVlVJaY4PlXLdQGm1t4AVppbmSLX33HXZ2sL5SMLFu18RfqcfHJ5R
p+Us5Mw9zKyxXgjuQdOut0arliBt7IQ6Oi0RW448YDev6tZ+PMTG9HeiPTKYZFxu
uZDSJrcOv62CrgsNRr8bkQCuGz45TC+PiYcCkGFU92t6bBYeWon4e0zSn2+NH52V
Vx0oakx2m3uKePykLx7joYGH0ejxmE7GcDUdpO4DGYS7DykejKbiQCs+d7vKMty2
6wBxzt89ziV+ekUQ7jE0lZNaMzByPevZ9Zq9mUnaPd3xTHdzRr8DpSpIi8h8WPIJ
WB1HGruK9CBXFGSeoITeWOaghRQpue4CeXhvBLBSjzjxY+LdEjBDubxuved7pOk3
q/AIUZM+cti0HN2cjFzfPJXdWvAe9tnEeWy5YieOJw7ktTDfOu86GuZAqz2D4SnD
mXuFelsoXoK0Y18FbeVMtnLfOQeltzkFsd0VomsHrm/gfeV3dsOa5MW2o6QOQM/8
jlhISiXFu56BE25tjzQ97p+SwGV+4XSlozN8u04PchQl9nkXQ2hA2sZBDqCLJZkT
qD0NLLLYJvcEpx3YZyYzV40ygz6mWsxgfcbSLbyjd4EOljRhK2DOhA+EvSpxB+WN
NyeO+KBxtQf8ENXkgqSD9Z/NiAmVGOhWve8T9PCXeTt6TRZkpFjLkvgunXKtrAAT
7GKvhfZJTQFyGTBEDWRrNnY5VbldIrjGS1pP/xRl0C1mwRNAQBeby8q7YB++QjYn
yGYLg112/chW/W0JCfFnGHCTqle5H4F8W28YCdCYaaMz6B7vdJgNPC8uevVORMPJ
Ahn6lSApK8bjfoEkiUNt7cy2VKrtO2kNbtW/AEZaflsKANmpolfJJQ/tMQT9v7Kd
GNdFcSL6uZEZ7UEokd6fJYo0p+najR2P+VUXplkoKGxgZUARvjKV6KEgTLhs3EGu
CiQSg+P2jM1dGA1yixOVnvD8KLK1R6t9S04uHGykEN1Asq6q1dKO974gIRHz4/ft
iIDsGCrGgzrOXrQiCy115TAsMrwAEAqYxOiBZ42yAhgTRbmLH1B4uZ0TjEZ0y2CL
1lbkcglz9xSaxwDS/KfBcrLcRiwRWnpoHg82CBg5mqxml7HtZ8XTS7qcnBK4XJSh
2IRh01BZd61jAp5we7b6IV9ly/6QWYM6EQXzk9v9Spw0E+kW1o+BxMGRyHPzja91
sPasR+WsvNCqt4tX5Tjj3lL1FTBwG/I4uT9bmiRGx6AMpH21eOMjDGkTLMa3Bt2h
ocywUJpHTqZrHmpR8ItnZm0Vsh3GzB8aKMM7xpAbK8maQqIzpnOrMRCzdpbXd8o1
dG5qmn5iIcvybLPpEF4j2FqbaAV6ZiDAG1Le/wcF5QKBg7fPFW47qhowPVifW3PT
g+iGqUudA70wTzq5jwlESPPSHiuFwXJWqQqrcMQPPZnqDSpllqKxOrf+mm/fNsQk
iP9wnl5tThKzgxns86OwMdeV04SHmOgybJjaV3rx97TtDYMR2AKF6VZc/IJn29m9
0+fyQkLcCcZr3o+2gEYhu4Is/imC21Yd4p/6LJ281CKOBou8Osk3gTO7+CLBWF/h
/B2JERoKt2NepCgyB4YGOyDPhedaq2NxrfchHJILpB4HxApPStUqzzp09qUC8IhK
GQfPi30tBx5xJNif+eAe6yLpn4rdmzCDqUokbbxhakGS4NtCRudahclS01x6J66v
jPPPqNvwb3xSrHf/GRfupDvtRVsiUcKiivF1KR1r+31JAwIczjTo0iPPOzHKr7v/
nraYeaevKBppgeh7vt+dQ/eXT5fVWtr45xZmyo1ukjdcX/lihUUSHlLTfpes100H
JFt+CZKa1wpuX8GBccD+C6F1hGNzjjcSKHrKoob/yCsDChsM7/2b+L3H4emokkI/
kL5TDxr6X1OHTK89FT5BDcpYPVH7CTbC76CWZcia/RJtfXMBFSoVeDEElVPMBAnv
vlbtcMpVLrOTHwGGcSzr/nncbocfriN1XsEB5+lwUXdRbUDjuxYPfd6qQjnvP8dd
PFDcoz5tFm/bFsRcYHoty3DqQWMVUStyMX1n5h+IXOAVHMQqWmgz55E0uRPDgN0z
ZtYfh9qn/GoIlJX1ygJDSBXtAOgqr6/WeECGw+0ugc2CiWofotgiJPwz201SReix
tIdd/lTvN1jWcOke0rBUkJ3IBQsMIXqVzetEjIIAycl88V0IOl5htKaLZoByZPeA
U6hvoTbmB8slMMm9ZUXwKjgPNyZ+IpzVT9dD/d+Ifg9xE7azK25K9dSndwSbwi9S
5p4JycR8a0/v1D1vcgphWwsajjL1u6BnLn1xUx/n8EQLA3IlPF0DNIS54xuYjdqR
Zfe623cQXtN67UgOvQH9DcLJpj4IPyCdZ8QYYx0+ZbCSm8UqtbrMiz5qCZO1N8mx
xroglwOY6Tec7vRzVVkfRQdTbnVT3QV5QX2YNVF529Xkbr8Ue/tXdgCqPg983EIh
htPN5JjL1JlMQ1rW01xrz+gRDjX1VcTgjbl3V+l1aJ8LWTPk0dd5qa2YPVxif8Bj
31lQNbanjATH35Rfda3398aSOjr10ikm7r3y2tbzBd4+aWYkMtSyy70baSEiJfLW
u1nveeue/Prq4+y57Zo2Q3/j6z3aPOq5YraYV4CF01GCs/dodYMrQeUAw1EtppOF
e1wZ6vu5tnQvBUY3PknbX+zEuwQzpPczanRGBXCIpgLQXUvUunS83rEHjpGvBqRl
S2zUgU2T6u+vmsTGCxtRzJnKskkRFtnUAfD03RCt4FzhJqMm7AEbed1k0Bu8IJSy
Yve4EGZPP2vq6/5UiF/OYlk9p9lqVawCgVgXpu/aVCrQJ4UQ+kL6Xj15nq+MOBtt
/QYY2zZhyGj45Rxjo7jTdo9y/o13VigWr3Jhxg7ZY8Dcx6tWlba+LWfvOVzkqd8P
YmEFCcUH1h8FGvT//Xb4zmpD+jPtGNORi48WrNc3L4EUTktZdHUOY9Hgxg8/GAZd
eWILin66bskMXtjoBFyiNdG6gapZ8kcc0qMiNNRqq6RIXIG0xHqonZpKEJlwdXDg
UrKTrshGNGQ9vBixJ7x59u2K++cSSltiov9a4vmSTKRaJ2z0vO290aFS9AldOgHJ
VrBpC5wCHqd+ypoqD40tdvfF9hvvsmapHEGyNDygv7Gbudm7zlnemBVwclBU8rEz
2OsrvEKV9vs/ia1bKfB2TH5Ta8ZB7IvLp5qAAg9PafrZqrR8IMiGmKAoXOermiWo
eOUHoFLqPWA4hxjtbgkxwVkmcC3pxr1RvSJZOk1JChENGKQ+WQ+bz9vyy3IlPsyn
36SGLbm95eEsqe+AAjpYNZH7SAiM/d2n4YAta+TQz8vp/AQBddJXN2CJmmkTohGv
Ko2e/SIGi5drmHHEtDTcxyuScvm8U8l/ro8ZSWSkMIKsYSEPnuwAcLkMWn35cV2s
gO6SwiyyEKWWgaJaCRpr+RSUJQp2XhsKIvxLLTZmzOupoTaUxWhbXNr8LK1ZBb23
fJfCPiD55rbn9DL72HH54pW1J9Nh/EwSGLZoRF1FXxEl/lUKfQmXoT2P1jAwuczJ
gnOF9JjFdyT70wEkqJ4Fz+/pX9Gl9wQPuSMcAV4N1UAfQTDoHdra8u8jQTE4ursC
lGuHozGV+VJdM2LSUW4qb8ghtc/zttB5NeoNG8JYilYSagBojUvF7GTlnCjid21D
ADrVEgrKo1ANypIoJz89CVl4AJpUHq4zFBzwoLybOxIWeKEN1lNJy7tXATRHHhns
eeEBMswbGHu30j+oKR0KOx44Sos98bMHyX1l8rWbNXCGUsW6CfCZSKdNjg1qL92C
i+GF6rt/Ys1mcdzPUcVI/o1TLDdVnB58qesJDYuognsEt23kyTwwmbCnK2zgx9qH
8wtWyoQQ1gLJU3gq9t8ZfGVTLGko8oIP+6CPEo6pyK1+KBHeKXwL//8ifzxupAzu
Ibc/V/oZW5qMlz1fm/OPktsummh/1KuX71rs83DqjxY1TRy3eY18fxwWPUi8sOxs
tSIRmYqfiE00HOrCl0pigDvG/NgxXnZ+NRM6NMnlUJOpqTetUbYkHS5BARBN4ch5
sKT0CSmf/TaVHBdb6OwvMlOUkbxsgHKe8hFc87Xjg95Flc8Hf3x6YJ6i1cgKPIRj
jS+LFTRlHV9cS4lYMmlGmLVrprax8cRxUnBeePinLgfFt8cUXowS8gKKnuhyWYwv
hBVXa1o9sG5NyBoXgPuWF2DFEAirlkA8nc5BSm09p9jIObclefhikeddk1DXvv5T
FSM5Tvi51sAfxLcH/DA90fJFrT+hEbo6sa+VD5oklf4zzOpFGTbKgO+ZTavNbXP0
TPbIFHP6APcZfNx8vpkCfAWv4c7Qvr3c5Z3rpiAXz7UkRR8vVX07A4iE3RrJw9RJ
yUFtWuUvVxAdTSXbxpKgfaEj96/jVnT7X5Evc9MiGF9gPsicWrSTnPx9Zq1C0LVJ
Z0YXmaaFWvu3ORbcoC+dsNSi67I9eRSax9ZA+TcIO1NSoeoveM+SMZfgDrlwH01A
8XJcJdXm/9qds10Icid4IElr1eYqr1S1oKjiEttLmNFI4m6yu2E3EGLerKaumjKT
lNwwQKfJCPNi46UHbLGbxMJZu4jeNUlZMXA+P5Qo5C0nuLgo8INopkEg7d339iHn
jCI5dI5BfQDUHgqO3gRs77KFFXLYCm8fX6kvfxe7rsTdEgThfnw5pFwgWx1aIZMS
7xUtBVzod/MJLEilLoDmF5uwzVP5YqqcAylqAJRF0vkcqfxScHEEqvneS6kovSOr
ZER1jKYkWNTMElrWsvbK64bXPrNJlhQ1uorj0kRrdVi8UZzkVxht0JAmaqF6psWm
EKu+M3y0wObi3filu0DX6WXrXKxTru9thzGyjIIIuHPFYB+D/lHn3Oc5eXegxREw
Y9ElHWV0snwaOAdO5KEgp11Y3eVL2xR1Nuys50zG8kx4kr5SmJklUvbr0hpppHJ9
ggtaW51gG4HGod6TIWe8RX+dkfAqdWoG655YmbfWUYY2Vvq4AnyxtzLRTg3fFQtL
1kjTGX/3KdrT9CbDLEAPSgSmUVgXGIYGDH1UF4a9L9ergAqUorL80UKDZj9M93QH
zqcQ2zTYwi3mHJ/hLP6ouEMoKwwDMi0301AFmoSDNfNYqXHODjdLmOl3ZlbozESL
af7CIEXQgkGY5GNcidzg45gbAI8FJ8V6thxOlPfWmO6WZiH2Hjn5GI8IWpQr5FcU
ZZ7595ljDiRkQA4BE2JqyMmXQN/F+Bq9wU227MqqcvFWXphrMEkWQwDJZhcQCkpR
LHC43azY3SrO/nF0VlGfb3OHie5TeNJd5JqeJx3xSCLopYW2fjsrsF/1VuBeOCLI
AYvpEtwaQ4uTY1rscImKxrZb+O/zpm7rBVHwQ7wJ0j+OAETFp+BT+/cewIG6i4eW
pc1a1zrtvG6q3mBCf97DDg7uFiof3WcvInt2LIbl5xxcQEW4JgC1S2VIt6j06Ktr
cE/o6j9U+2/fL58dHlFAzGIK3sUaQCx9bcUBjSW8Rvrl0HT2c3/moTtSQbTqpT8v
0F01QFWOXS/Isp2ng99qSt+DhKnVQAEEG/ZjPVK5eFnBdWunN1YB/rUg71Mp5lN9
i/NH/BN53LK1srxmTV0f/s5itzUCo4qrULzm+B1WlqlSI+T01UPmO0EJdkM+Kx1K
r0R/SFGFw6qCvMztmDunyia56MdHkvPG2gmjGaig5mQnXkL7zU0K4RXfRtBkiON/
7OsFYT4d/cPN/ni8Ve8w4NiCOnSpZ/8OF/B0DnsiGrss4Kpaad9SPMzfAejm1+n5
q9Ix2iptLJuS/pw5EfkOGpoeie4F052+C734MMTGlq5xZoD2+s4tRK05JN5aqrih
qegWeb3csxaAG7cOlxOEh49Q1ngWN89QYJBpf791iJEFaZLfYkuS7O+XK5ZTu2gp
JP4dEFiU08lQXqMbFsYM87xU5IoPEYww2ov3cmBLZrr8iPoSJm0Uk/wHplXY1RHT
A5mX4O3YOfH6LWOSCHJNXN6Mc8YzMTCOk2evAp4OGzXOC5OBWtfGUDyvfrKozMI/
QfG4hja3ySQQhFblxi55y4XJdvMjzO1E24m80VL5yBrGK6evW3v2rDydyGbisV9V
WF2jjN1B73anjC87VEa0hNfiqlrk4jDh+Fh4PpHRkkcW1/dJimCLDHTA0qdon7aP
DC0FTveR4JPSqS0esyl9zIjVWP/ApMoUqupiq9Sg5mSfERHytFKOpWUk2pvA+R9G
8TP9+inCp7exG/bkDh6kfWi4pV5lXtl6cN56e0W04xz6xKorqbm6tOp5DRZsjdzu
bjTeXuBpEEfle9P0QPjp+doTk1f3ib3JnAE7k5uQzZI1W86Hqw+Akkl92+hw4xcz
iL4dIN5hfLmTA98Nqo3a4rdnJbByOdTBetUTRZQoPzxdDrrK07FMk3PfGj5C71Er
wFvYZtFhPd8JfsoDxEW1kLvtbPatZ7KSRePqjsO5vBv0DAEfmQDS2lZJA7goICEp
k4oqogkpCEAedaJenARnH5nDzMkJvwAWToeKTI7cTA6hco33bKGnZi+8238P76Ot
RHBBXOAdscvP0Gu7GBJY4mbXg99ArJOF8oVKdwCjzO8iADwzzuSSvwbS2WZ56bdh
IDqrS5lj3OeY8n29LEmDXDMvxpgjB9n3AnnMump9DsnwuVvvWYoTPOtkQdysetb/
gMeLoQLJJvBwgR4b8cqel9tjsSUQqOf7piMoiUXqA4RDST6yqISJRCn4gCxXFKYJ
tUROx1VTHLWD2XXNyR8Kza8BJn/2ykg381XUTGia2tbBqBhN3TPU5/Gt/gw8qkz0
Mnk1QwDLNqf6FprWx6sU1QVW2oJo+pDFahNVNcIPtUo6BvUTDZuqIcTZtpKaeYBW
CtM5O/d3nPNNakPeLApmTg4Ok++8EcvQmxQL/bIo33c14l3AzAbbyNvPn9gEjJU1
HMDcCgerpfcaE+QvelsEtSzcBDSspubJ/7xx4xzVdEghCugXH9XAcjdopWXWmOsx
LwOK9oHI8V3DqEI7ldODRQcciXa8prboiZMuIaif9Mret8Ib8J/iB5iBuJLUxJEJ
yqNfWpVZ2KGLDKX/L11HKXBhIxjAxprvPZt5Cb+GOgsgXKxuH8SjvGRdSDNvAhKt
b3L+C0NC32zjfcXU57QR0AxNK8wY4vBv4l6aqS1nnQsoBlvAiVUBvZGDL2RQqr1s
7lrPaNlAvMgxIFsigD8oEsRx0xuOjf0HgxHzgkdVohvol4kbuBOX+CTzFAICx71C
zcirKS9JkM07vdbZKxBHp6H4iX4ZQauARRiMIqPcqxAaaWiBwKO/y22tatY+f0uR
44e4HxYSB4tla1Mq2BCivpodyna9/UmUGQZxqVi41020qhTD9SvDIH3ge1ARnwm1
GDrHtkbxQz0LmbPTy3LPcL11tNWQ7UGdSaZbHX2UUw62lf4var0s7Rw2bEkyAx3v
Z6MRDKQitPUYEUyspgWu99HtdptcW3Q+g+SoKMvD0j4u4TxxB88uSlsnzPtqTN9r
zbolVL479MfcaFtzC4BJhpbgcscYhhheZWcut95AGDDeZoNOMEuvEarPUXlet3Vk
oUD/0XZ1nhFsK43Gjn2x4Aprbz3DZDjOsR9iWNyrIkGJp40DqjDj8N/jmejwxkW9
1QCaYN4Px2sfXrVE927HNeFtEp3+ofNi6sffaIUcHmrPt89qu7EoKbnMJhblPfBX
zQSmSAdyJ7/hCDkZFU1BQ2hlyHI6imAQUvxq7QFGswhgA44WQ5wzaPp3RfoAMvSC
+Y859hbZmbwhOaR1Tby+DhABcNhE96ehNqo3oSGUpEA8G53rlugcrNntsJ34ren7
/aqcZ7dFpdFbHYJq6cgZqjAjcGdl3kV8gAsPcZQTxDG03slV1nxNPJApH9lH2WZL
XtGCk3AZDJBGEUKyFpShSTKQdiqUTXBZNaHCoUGxvgviqmkx4eHNGiu9YgPIczZH
NI8dhzgFShDxLpHDg5mpoxzemVr6knFzz9Fqgebrx7wDhBRpo6fpP2X/E0Q+A5fh
rZek1thLg+qk7wywcR2BaHulfWNmJ5PJfCnkwNyZXZEb3mqVBOkE15vdhRy+7RU6
QUQcGRGam9GK0B7rpH7wB0xOh+ql8RUdlwPZTfvq2m8E3OO09Ih3W4JE9hO8EiT6
l4WjEa4fEdICmcdg7c01EbLj5mOP6e4XpL87ZcXJ7Zb6s3DQcPBBBEyDIsyz6cq+
cupsxizAYsVqS1VKot1JF/XNf5u2Nv65l5QeqR2AHrRJ1CqOcGeSFps4GkhSuD4S
1pNif7BYQxBbJfENvFyf3oOdcC0TqIEbp8gumRWXOtbssEjdmaWvQ/Any+xW4EpZ
fXziaSMwMkJdVphQ9IdRTTmPdDrscnFuYhEWj1ewk5/DiJsadvshORS61kM4yJ3A
6sdBmMjbVMKfsM3mUgWjt6+QRCa7l1npjL2YUwvE79hVXHvoiKlndWI7MFC8s2ph
f+Dm4S/6oUdySZbq2zKClyioa/c/c27C900pEWsDBHv3E4uLzJbM0Fi7X9CcDpo7
S88NzkBtFCswcUvDSeclssJg/6ERJpbynT2GalQgRpyvjdo7+8bwkRwFl+p97Ejx
kllh+8onvAZCJ7VOmXMkTSvj2myNdzFElPHLToJx+rEjN6wZqt4xiZVOTT6dFh8Z
erGjb/quBbgJDH55SqJIbrY5dNJyst/eqUr3ZIES3eDazHMTNqV8aE4Nf9KgKD0U
ZlnCGifN9VfrQObQkkMfHLGG07VHhoQgt2DjcdtC5IIZ4BUKwkd2NfVnaj9qL12t
bhhhZRqHtKcnR+2AL1+1eHs6r+uKhOv8TU9stScrKTJrQnZlBbUWg/kUunw2jwzk
XDStzJPCv9ArVkf9ZV25XDk1nMgGi+vuJEWbLnU3vJVXOxAlbfb/cOU6ulKkil6L
QkdDrGl6uigLIzd+ZwhQrshQcGjR7vGoqsBaBDNbzmDZa1cmPYjsPaVVQI2q3Y8m
ei0t6paTIeLqv8nj3RwL7b9y3LFJJ1WeglsW8qJ73o8dXCegRAm3MaTD/XvjtoiG
dlH4zyUPDvXmLXt5b08H6CH0D7EQMHkP9HYRo66eQEXcQYgF+yaDGqY7jjNH10Ec
CHUqUtdda5dhYtGbJiHClpnUK/GsdTqPMYOFIz8QUWp9032iY0PPDakksLWNgWM9
/y6ZdIlp5aU5X5bwkyhJLPfzJ73oUaRz78yZ5ZTEkr9GqtDSqsUc0S6vaFgNDG4L
fPTDmLFVgBnMycSF0Mx/B46IoPRA3mae4mLWGzL86GkkBmjDL4S/N8gCeCMh/AdF
uN693pT7e8pFBsokMaf73wwgvV9WJiti7S6PJHdnmrCXDyDTgFBmEpQQV2Wme9zI
hCWUIUgCLvq4uDq/o4ogKxS4Lox4yX7HqEsmbFOTdQP5Xn+Y9IQhsErGZR9JGEuq
3ortVrmpTzlwdF1o96Lf1d6VwEY3dCQPSbf+ElTyv58G5cmqShcalYwJgmM+3zqR
7vcgy+9kfUUKngoEtZgRbuHr5wrnVn9EsKs7GodprIlF2W8o1bmR4UNRNmXNO7eD
MxXEoIYxjsDZP/agYINNlTRQ11q4Yw9UKH48iYkQ/chaUiABvuivrOnCqVQNKGWr
80l878z6+/f0ORZrwn8iHJLDMSJree1Tu/ghByvmw0N/yjPcYe4V03yE15OhsaDb
xauEar4D8WClnGxxpn/FMspMr4qF/dwxMpk4ZB/7MNGpTFfyCkj6iANvT40VAEJr
0tDRmUs8Rf6s7yi5bpR2ZArcNrcw3RMpnaPbkA8/WC4GBKmulIcEMzO1jJWkNDpp
MmtCt1TZZufj2bC90kSgQKombE69wKHRPNtwzn11lldJxANeV1t0EL0AonTIhjth
C1exrbsUQRYnkiHHDiAOWJFQ9FofUaSvFZ0MZoQkfMH46gHn5/AVRQE5Nu6EY5r8
ZCqhOj61TbBfRR8WASBNoW69xsQnpIkEdfXkyPMf6S3KLLyrn4WTlsB2mKEOwbLj
qgh7SCHnK6j25xS/x8q3lAolixmGMa8czwlstXAiM9/mqhOb4UDSzNScmHG/gEEm
4k3E0+z2kodwK6n+xbJOK+bbeeNpw8CojYBvAoddqIkBYJ57Xt4Yjj7pvSNwXdtz
VzEIi5nvt5ZLqEjV4dmXmtSWI0j1Sk9c1+/81PNpHe9j++C9OyRLNu3Z5AYn38k+
NGBsJZ/fbdSstvauP6Il3Hhz1hcwKfxgh9IjFzDcXIK1sWGGgg7sZzdQ2VxReORD
1MAD17ABEjEle5KX2lFGD2nX7Uc2APE65JWvnSm/3WokccFK48F3MN5IPGSXIpjM
ZFhPd4P6EDGoEZplSFWFaA==
`pragma protect end_protected
